ex2.vh line1
ex2.vh line2
