included line 1
included line 2
//>  incl_file  "corpus/ex2.vh" 
included line 4
included line 5
